`timescale  1ns/1ps

`define     DATA_WID    10
`define     WN_WID      10
`define     ACC_LEN     8

// `define     FFT_LEN     8
// `define     LOG2_FFT_LEN 3

// `define     FFT_LEN     16
// `define     LOG2_FFT_LEN 4

// `define     FFT_LEN     32
// `define     LOG2_FFT_LEN 5

`define     FFT_LEN     64
`define     LOG2_FFT_LEN 6

`define     STG_WID     4

`define     WN_LEN      (`FFT_LEN/2)



//------------------------------------------------------------------------------
    //
    //  Filename       : fft_core8.v
    //  Author         : LiuXun
    //  Created        : 2020-08-02
    //  Description    : FFT core. 8 points FFT based on core2
    //                   
//------------------------------------------------------------------------------

module fft_core8(
    fft_i,
    wn_i,
    fft_o
  );

//*** PARAMETER ****************************************************************


//*** INPUT/OUTPUT *************************************************************
  

//*** WIRE/REG *****************************************************************


//*** MAIN BODY ****************************************************************


endmodule
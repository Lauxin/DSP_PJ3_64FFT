`timescale  1ns/1ps

`define     DATA_WD         (DATA_RE_WD+DATA_IM_WD)
  `define     DATA_RE_WD      10
  `define     DATA_IM_WD      10
`define     CFG_WN_WD       10
`define     DATA_FRA_WD       8
  
`define     SIZE_FFT        64
`define     LOG2_SIZE_FFT   6
`define     SIZE_GRP        8



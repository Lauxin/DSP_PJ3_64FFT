`timescale  1ns/1ps

`define     DATA_FFT_WD           10      // (DATA_RE_WD+DATA_IM_WD)
  `define     DATA_FFT_RE_WD        10
  `define     DATA_FFT_IM_WD        10
`define     CFG_WN_WD             10      // (CFG_WN_RE_WD+CFG_WN_IM_WD)
  `define     CFG_WN_RE_WD          10
  `define     CFG_WN_IM_WD          10
`define     DATA_FRA_WD           8

`define     SIZE_FFT              64
`define     LOG2_SIZE_FFT         6
`define     SIZE_GRP              8


